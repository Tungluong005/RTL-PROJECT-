`timescale 1ns / 1ps


module NOT_GATE(
  a,
  y
);
  input a;
  output y;
  wire a;
  wire y;
  assign y = ~a;
  endmodule