`timescale 1ns / 1ps

module NAND_testbench();
  reg a, b;
  wire y;
 // khoi tao DUT
 NAND_gate dut(
  .a(a),
  .b(b),
  .y(y)
 );
  // Khoi tao Stimulus
  initial begin
  #0;  a = 0; b = 0;
  #10; a = 0;  b = 1;
  #10; a = 1;  b = 0;
  #10; a = 1;  b= 1;
  #10; $finish;
  end
  // Khoi tao monitor
  initial
    $monitor("a = %b, b = %b, y = %b",a ,b ,y);
  endmodule