`timescale 1ns / 1ps


module And_gate(
   x,
   y,
   z,
);
  input x;
  input y;
  output z;
  wire x;
  wire y;
  wire z;
  assign z = x & y;
  endmodule